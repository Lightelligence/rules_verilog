package apb_pkg;

   localparam ADDR_WIDTH=12;
   
endpackage : apb_pkg
