package dpi_pkg;

   import "DPI-C" function void echo_hello();
   
endpackage : dpi_pkg
