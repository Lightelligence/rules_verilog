module apb;

   initial begin
      $display("apb addr_width:", apb_pkg::ADDR_WIDTH);
   end
   
endmodule : apb
