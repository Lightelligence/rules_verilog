module unit_test_top ();

   apb u_apb();

endmodule : unit_test_top
