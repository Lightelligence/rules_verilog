module apb;

   initial begin
      $display("apb");
   end
   
endmodule : apb
